`timescale 1ns /1ps


module ALU(A,
           B,
           Result,
           ALUControl,
           OverFlow,
           Carry,
           Zero,
           Negative);

           input [31:0]A,B;//Declaring inputs
           
           input [2:0]ALUControl;//Total 8 combinations(or 8 operations)
           
           output Carry,OverFlow,Zero,Negative; //Declaring these for checking the overflow condition, as well as zero carry negative flag.
           
           output [31:0]Result; // To store result

           wire Cout;
           wire [31:0]Sum;

           assign {Cout,Sum} = (ALUControl[0] == 1'b0) ? A + B :(A + ((~B)+1)) ; // Subtracting using 2's Complement and using Ternary operator to generate MUX           
           
           assign Result = (ALUControl == 3'b000) ? Sum :
                    (ALUControl == 3'b001) ? Sum :
                    (ALUControl == 3'b010) ? A & B :
                    (ALUControl == 3'b011) ? A | B :
                    (ALUControl == 3'b101) ? {{31{1'b0}},(Sum[31])} : {32{1'b0}};
    
           assign OverFlow = ((Sum[31] ^ A[31]) & 
                      (~(ALUControl[0] ^ B[31] ^ A[31])) &
                      (~ALUControl[1]));
           assign Carry = ((~ALUControl[1]) & Cout);
           assign Zero = &(~Result);
           assign Negative = Result[31];

endmodule
